module spi_peripheral (
    input  wire       clk,      
    input  wire       rst_n,   
    input  wire       nCS,   
    input  wire       COPI,  
    input  wire       SCLK,  

    output reg  [7:0] en_reg_out_7_0,
    output reg  [7:0] en_reg_out_15_8,
    output reg  [7:0] en_reg_pwm_7_0,
    output reg  [7:0] en_reg_pwm_15_8,
    output reg  [7:0] pwm_duty_cycle,
    output reg  [7:0] uo_out       // <- exposed for testbench
);

    // 2-stage input synchronizers
    reg nCS_sync1, nCS_sync2;
    reg SCLK_sync1, SCLK_sync2;
    reg COPI_sync1, COPI_sync2;

    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            nCS_sync1 <= 1'b1; nCS_sync2 <= 1'b1;
            SCLK_sync1 <= 1'b0; SCLK_sync2 <= 1'b0;
            COPI_sync1 <= 1'b0; COPI_sync2 <= 1'b0;
        end else begin
            nCS_sync1 <= nCS; nCS_sync2 <= nCS_sync1;
            SCLK_sync1 <= SCLK; SCLK_sync2 <= SCLK_sync1;
            COPI_sync1 <= COPI; COPI_sync2 <= COPI_sync1;
        end
    end

    // edge detection
    reg SCLK_prev;
    wire SCLK_rising = (SCLK_sync2 == 1'b1) && (SCLK_prev == 1'b0);
    always @(posedge clk or negedge rst_n) SCLK_prev <= (rst_n) ? SCLK_sync2 : 1'b0;

    reg nCS_prev;
    wire nCS_negedge = (nCS_sync2 == 1'b0) && (nCS_prev == 1'b1);
    wire nCS_posedge = (nCS_sync2 == 1'b1) && (nCS_prev == 1'b0);
    always @(posedge clk or negedge rst_n) nCS_prev <= (rst_n) ? nCS_sync2 : 1'b1;

    // SPI transaction tracking
    reg [15:0] shift_register;
    reg [4:0]  bit_count;
    reg        frame_valid;
    reg        transaction_processed;

    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            shift_register <= 16'd0;
            bit_count <= 5'd0;
            frame_valid <= 1'b0;
            transaction_processed <= 1'b0;
        end else begin
            // start of transaction
            if(nCS_negedge) begin
                bit_count <= 5'd0;
                frame_valid <= 1'b0;
            end

            // shift in bits on SCLK rising edge
            if(nCS_sync2 == 1'b0 && SCLK_rising) begin
                shift_register <= {shift_register[14:0], COPI_sync2};
                bit_count <= bit_count + 5'd1;
            end

            // end of transaction
            if(nCS_posedge) begin
                if(bit_count == 5'd16) frame_valid <= 1'b1;
                bit_count <= 5'd0;
            end
        end
    end

    // commit to output registers
    localparam MAX_ADDRESS = 7'd4;
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            en_reg_out_7_0   <= 8'h00;
            en_reg_out_15_8  <= 8'h00;
            en_reg_pwm_7_0   <= 8'h00;
            en_reg_pwm_15_8  <= 8'h00;
            pwm_duty_cycle   <= 8'h00;
            uo_out           <= 8'h00;
        end else if(frame_valid && !transaction_processed) begin
            if(shift_register[15] == 1'b1 && shift_register[14:8] <= MAX_ADDRESS) begin
                case(shift_register[14:8])
                    7'd0: en_reg_out_7_0  <= shift_register[7:0];
                    7'd1: en_reg_out_15_8 <= shift_register[7:0];
                    7'd2: en_reg_pwm_7_0  <= shift_register[7:0];
                    7'd3: en_reg_pwm_15_8 <= shift_register[7:0];
                    7'd4: pwm_duty_cycle  <= shift_register[7:0];
                    default: ;
                endcase
            end
            transaction_processed <= 1'b1;
        end else if(transaction_processed) begin
            transaction_processed <= 1'b0;
        end

        uo_out <= en_reg_out_7_0;
    end

endmodule
